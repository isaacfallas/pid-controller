// Code your design here
`include "PID.v"
`include "16x16bit_multiplier_pipelined.v"
`include "booth.v"
`include "CLA_fixed.v"

interface intf_wb (input clk);
  
  logic TAG_s2m;
  logic TAG_m2s;
  logic ERR_s2m;
  logic RTY_s2m;
  logic SEL_m2s;
  
endinterface

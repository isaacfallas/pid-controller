// Code your testbench here
// or browse Examples
`include "wb_master.v"
`include "interface_PID.sv"
`include "interface_wb.sv"
`include "PID_tb.v"